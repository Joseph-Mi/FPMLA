module main (
	input CLOCK_50,
	
);

	
endmodule 